//------------------------------------------------------------------
// Project  : EDB HDL WS2021 - Fifth Assignment
// Purpose  : Implement a testbench for an UART receive (uart_rx)
// Author   : SteDun
// Version  : V1.0 2021-12-10
//------------------------------------------------------------------

module tb_uart_rx
();

// (1) DUT wiring
// (2) DUT instance
// (3) DUT stimulation

endmodule