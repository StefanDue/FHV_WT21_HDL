// ------------------------------------------
// Project:     EDB HDL WT2021
// Purpose:     Implement a testbench for a finite state machine door
// Author:      SteDun
// Version:     V1.0 2021-12-10
// ------------------------------------------